
module hello(input clk);

initial
begin: proc_he
        $display("hello 1");                                                                                           
        $display("hello2");			                                                                             
end

endmodule
